module input(